//!The module is used to simulate a mmu module ,**only for testing**.
//!              The internal implementation is not the same as the real mmu module.
//!              it will use fifo to store the 4K page addr, so the address always
//!              be the 4K aligned.