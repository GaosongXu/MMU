//!connect to the fifo, and filter the invalid requests
//!do a dispatcher and control the switch between the alloc and free mode
//it will maintain a fsm to control the dispatch logic
module dispatcher(

);

endmodule